//--- Parameters for register addresses
localparam   SNVS_ADDR_HPLR     = 12'h000;
localparam   SNVS_ADDR_HPCOMR   = 12'h004;
localparam   SNVS_ADDR_HPCR     = 12'h008;
localparam   SNVS_ADDR_HPSICR   = 12'h00C;
localparam   SNVS_ADDR_HPSVCR   = 12'h010;
localparam   SNVS_ADDR_HPSR     = 12'h014;
localparam   SNVS_ADDR_HPSVSR   = 12'h018;
localparam   SNVS_ADDR_HPHACIVR = 12'h01C;
localparam   SNVS_ADDR_HPHACR   = 12'h020;
localparam   SNVS_ADDR_HPRTCMR  = 12'h024;
localparam   SNVS_ADDR_HPRTCLR  = 12'h028;
localparam   SNVS_ADDR_HPTAMR   = 12'h02C;
localparam   SNVS_ADDR_HPTALR   = 12'h030;
localparam   SNVS_ADDR_LPLR     = 12'h034;
localparam   SNVS_ADDR_LPCR     = 12'h038;
localparam   SNVS_ADDR_LPMKCR   = 12'h03C;
localparam   SNVS_ADDR_LPSVCR   = 12'h040;
localparam   SNVS_ADDR_LPTGFCR  = 12'h044;
localparam   SNVS_ADDR_LPTDCR   = 12'h048;
localparam   SNVS_ADDR_LPSR     = 12'h04C;
localparam   SNVS_ADDR_LPSRTCMR = 12'h050;
localparam   SNVS_ADDR_LPSRTCLR = 12'h054;
localparam   SNVS_ADDR_LPTAR    = 12'h058;
localparam   SNVS_ADDR_LPSMCMR  = 12'h05C;
localparam   SNVS_ADDR_LPSMCLR  = 12'h060;
localparam   SNVS_ADDR_LPPGDR   = 12'h064;
localparam   SNVS_ADDR_LPGPR    = 12'h068;
localparam   SNVS_ADDR_LPZMKR0  = 12'h06C;
localparam   SNVS_ADDR_LPZMKR1  = 12'h070;
localparam   SNVS_ADDR_LPZMKR2  = 12'h074;
localparam   SNVS_ADDR_LPZMKR3  = 12'h078;
localparam   SNVS_ADDR_LPZMKR4  = 12'h07C;
localparam   SNVS_ADDR_LPZMKR5  = 12'h080;
localparam   SNVS_ADDR_LPZMKR6  = 12'h084;
localparam   SNVS_ADDR_LPZMKR7  = 12'h088;
localparam   SNVS_ADDR_LPGPR0   = 12'h090;
localparam   SNVS_ADDR_LPGPR1   = 12'h094;
localparam   SNVS_ADDR_LPGPR2   = 12'h098;
localparam   SNVS_ADDR_LPGPR3   = 12'h09C;
localparam   SNVS_ADDR_LPTDCR1  = 12'h0A0;
localparam   SNVS_ADDR_LPTDSR   = 12'h0A4;
localparam   SNVS_ADDR_LPTGFCR1 = 12'h0A8;
localparam   SNVS_ADDR_LPTGFCR2 = 12'h0AC;
localparam   SNVS_ADDR_LPAT1    = 12'h0C0;
localparam   SNVS_ADDR_LPAT2    = 12'h0C4;
localparam   SNVS_ADDR_LPAT3    = 12'h0C8;
localparam   SNVS_ADDR_LPAT4    = 12'h0CC;
localparam   SNVS_ADDR_LPAT5    = 12'h0D0;
localparam   SNVS_ADDR_LPATCTL  = 12'h0E0;
localparam   SNVS_ADDR_LPATCLKCTL  = 12'h0E4;
localparam   SNVS_ADDR_LPATRC1R = 12'h0E8;
localparam   SNVS_ADDR_LPATRC2R = 12'h0EC;
localparam   SNVS_ADDR_HPVIDR1  = 12'hBF8;
localparam   SNVS_ADDR_HPVIDR2  = 12'hBFC;

//--- Parameters for the register selections - used by the address decoder
localparam   SNVS_REG_HPLR       = 0;
localparam   SNVS_REG_HPCOMR     = SNVS_REG_HPLR     + 1;
localparam   SNVS_REG_HPCR       = SNVS_REG_HPCOMR   + 1;
localparam   SNVS_REG_HPSICR     = SNVS_REG_HPCR     + 1;
localparam   SNVS_REG_HPSVCR     = SNVS_REG_HPSICR   + 1;
localparam   SNVS_REG_HPSR       = SNVS_REG_HPSVCR   + 1;
localparam   SNVS_REG_HPSVSR     = SNVS_REG_HPSR     + 1;
localparam   SNVS_REG_HPHACIVR   = SNVS_REG_HPSVSR   + 1;
localparam   SNVS_REG_HPHACR     = SNVS_REG_HPHACIVR + 1;
localparam   SNVS_REG_HPRTCMR    = SNVS_REG_HPHACR   + 1;
localparam   SNVS_REG_HPRTCLR    = SNVS_REG_HPRTCMR  + 1;
localparam   SNVS_REG_HPTAMR     = SNVS_REG_HPRTCLR  + 1;
localparam   SNVS_REG_HPTALR     = SNVS_REG_HPTAMR   + 1;
localparam   SNVS_REG_LPLR       = SNVS_REG_HPTALR   + 1;
localparam   SNVS_REG_LPCR       = SNVS_REG_LPLR     + 1;
localparam   SNVS_REG_LPMKCR     = SNVS_REG_LPCR     + 1;
localparam   SNVS_REG_LPSVCR     = SNVS_REG_LPMKCR   + 1;
localparam   SNVS_REG_LPSR       = SNVS_REG_LPSVCR   + 1;
localparam   SNVS_REG_LPTGFCR    = SNVS_REG_LPSR     + 1;
localparam   SNVS_REG_LPTDCR     = SNVS_REG_LPTGFCR  + 1;
localparam   SNVS_REG_LPSRTCMR   = SNVS_REG_LPTDCR   + 1;
localparam   SNVS_REG_LPSRTCLR   = SNVS_REG_LPSRTCMR + 1;
localparam   SNVS_REG_LPTAR      = SNVS_REG_LPSRTCLR + 1;
localparam   SNVS_REG_LPSMCMR    = SNVS_REG_LPTAR    + 1;
localparam   SNVS_REG_LPSMCLR    = SNVS_REG_LPSMCMR  + 1;
localparam   SNVS_REG_LPPGDR     = SNVS_REG_LPSMCLR  + 1;
localparam   SNVS_REG_LPGPR      = SNVS_REG_LPPGDR   + 1;
localparam   SNVS_REG_LPZMKR0    = SNVS_REG_LPGPR    + 1;
localparam   SNVS_REG_LPZMKR1    = SNVS_REG_LPZMKR0  + 1;
localparam   SNVS_REG_LPZMKR2    = SNVS_REG_LPZMKR1  + 1;
localparam   SNVS_REG_LPZMKR3    = SNVS_REG_LPZMKR2  + 1;
localparam   SNVS_REG_LPZMKR4    = SNVS_REG_LPZMKR3  + 1;
localparam   SNVS_REG_LPZMKR5    = SNVS_REG_LPZMKR4  + 1;
localparam   SNVS_REG_LPZMKR6    = SNVS_REG_LPZMKR5  + 1;
localparam   SNVS_REG_LPZMKR7    = SNVS_REG_LPZMKR6  + 1;
localparam   SNVS_REG_HPVIDR1    = SNVS_REG_LPZMKR7  + 1;
localparam   SNVS_REG_HPVIDR2    = SNVS_REG_HPVIDR1  + 1;
localparam   SNVS_REG_LPGPR0     = SNVS_REG_HPVIDR2  + 1;
localparam   SNVS_REG_LPGPR1     = SNVS_REG_LPGPR0   + 1;
localparam   SNVS_REG_LPGPR2     = SNVS_REG_LPGPR1   + 1;
localparam   SNVS_REG_LPGPR3     = SNVS_REG_LPGPR2   + 1;
localparam   SNVS_REG_LPTDCR1    = SNVS_REG_LPGPR3   + 1;
localparam   SNVS_REG_LPTDSR     = SNVS_REG_LPTDCR1  + 1;
localparam   SNVS_REG_LPTGFCR1   = SNVS_REG_LPTDSR   + 1;
localparam   SNVS_REG_LPTGFCR2   = SNVS_REG_LPTGFCR1 + 1;
localparam   SNVS_REG_LPAT1      = SNVS_REG_LPTGFCR2 + 1;
localparam   SNVS_REG_LPAT2      = SNVS_REG_LPAT1    + 1;
localparam   SNVS_REG_LPAT3      = SNVS_REG_LPAT2    + 1;
localparam   SNVS_REG_LPAT4      = SNVS_REG_LPAT3    + 1;
localparam   SNVS_REG_LPAT5      = SNVS_REG_LPAT4    + 1;
localparam   SNVS_REG_LPATCTL    = SNVS_REG_LPAT5    + 1;
localparam   SNVS_REG_LPATCLKCTL = SNVS_REG_LPATCTL  + 1;
localparam   SNVS_REG_LPATRC1R   = SNVS_REG_LPATCLKCTL  + 1;
localparam   SNVS_REG_LPATRC2R   = SNVS_REG_LPATRC1R + 1;
localparam   SNVS_REG_NUMBER     = SNVS_REG_LPATRC2R + 1;

// System wide defines
localparam SNVS_DATA_WIDTH = 32;
localparam [SNVS_DATA_WIDTH-1:0] SNVS_DATA_WIDTH_ZERO = 0;
localparam SNVS_DATA_DWIDTH = SNVS_DATA_WIDTH*2;

localparam SNVS_ADDR_WIDTH = 12;
localparam [SNVS_ADDR_WIDTH-1:0] SNVS_ADDR_WIDTH_ZERO = 0;

localparam SNVS_HACC_WIDTH = 32;
localparam [SNVS_HACC_WIDTH-1:0] SNVS_HACC_WIDTH_ONE = 1;

localparam SNVS_ZMK_WIDTH = 256;

